module	ARM_Pipelined_PC_Logic
	(input logic);


endmodule


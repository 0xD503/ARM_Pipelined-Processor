module ARM_Pipelined_InstructionDecoder
	(input logic);


endmodule


module ConditionUnit
	(input logic		i_Flag_Write_Execute, i_Cond_Execute,
	input logic[3:0]	i_Flags_Execute,

	output logic[3:0]	o_Flags,
	output logic		o_CondEx_Execute);



endmodule


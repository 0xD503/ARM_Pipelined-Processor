module ARM_Pipelined_ALUDecoder
	(input logic	);

endmodule


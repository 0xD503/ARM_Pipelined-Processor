module ARM_Pipelined_Controller
	#(parameter	BusWidth	= 32)
	(input logic			

	//	
	);



endmodule



module ARM_Pipelined_Decoder
	(input logic		

	//	
	);



endmodule

module ARM_Pipelined_MainFSM
	(input logic		);


endmodule

module ARM_Pipelined_ALUDecoder
	(input logic	);

endmodule

module ARM_Pipelined_InstructionDecoder
	(input logic);


endmodule

module	ARM_Pipelined_PC_Logic
	(input logic);


endmodule



module ARM_Pipelined_ConditionalLogic
	(input logic		);


endmodule

module ARM_Pipelined_ConditionCheck
	(input logic);


endmodule


module ARM_Pipelined_HazardUnit
	(input logic);

endmodule


module ARM_Pipelined_ConditionalLogic
	(input logic		);


endmodule


module ARM_Pipelined_Datapath
	#(parameter	BusWidth	= 32)
	(input logic			);


endmodule


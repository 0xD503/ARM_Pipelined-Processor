module ARM_Pipelined_ConditionCheck
	(input logic);


endmodule


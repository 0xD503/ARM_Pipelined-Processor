module ARM_Pipelined_Decoder
	(input logic		

	//	
	);



endmodule


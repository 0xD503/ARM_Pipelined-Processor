module ARM_Memory
	();

endmodule


module ARM_Pipelined_CPU
	#(parameter	BusWidth	= 32)
	(input logic					i_CLK, i_NRESET,);


endmodule

module ARM_Pipelined_Controller
	#(parameter	BusWidth	= 32)
	(input logic			

	//	
	);



endmodule




module ARM_Pipelined_MainFSM
	(input logic		);


endmodule

